* C:\Users\CS Net Games\Desktop\4th 2ndSem\Electro lab\circuits\Prelab6N31.scv

* Schematics Version 9.1 - Web Update 1
* Sun Mar 24 05:11:18 2024



** Analysis setup **
.tran 0ns 2ms 0 10u
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Prelab6N31.net"
.INC "Prelab6N31.als"


.probe


.END
