* C:\Users\CS Net Games\Desktop\4th 2ndSem\Electro lab\circuits\CMNEmitte1r.sch

* Schematics Version 9.1 - Web Update 1
* Tue Apr 02 16:26:22 2024



** Analysis setup **
.tran 0ns 50ms 0 11u
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "CMNEmitte1r.net"
.INC "CMNEmitte1r.als"


.probe


.END
