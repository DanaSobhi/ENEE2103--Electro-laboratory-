* C:\Users\CS Net Games\Desktop\4th 2ndSem\Electro lab\circuits\CBase.sch

* Schematics Version 9.1 - Web Update 1
* Sat Mar 30 17:46:20 2024



** Analysis setup **
.tran 0ns 50ms 0 15u
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "CBase.net"
.INC "CBase.als"


.probe


.END
