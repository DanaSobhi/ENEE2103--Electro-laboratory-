* C:\Users\CS Net Games\Desktop\4th 2ndSem\Electro lab\circuits\Schematic5Prelab2.sch

* Schematics Version 9.1 - Web Update 1
* Sat Mar 02 23:01:02 2024



** Analysis setup **
.ac LIN 101 10 1.00K
.tran 0ms 100ms 0 10u
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic5Prelab2.net"
.INC "Schematic5Prelab2.als"


.probe


.END
