* C:\Users\CS Net Games\Desktop\4th 2ndSem\Electro lab\circuits\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Sat Mar 02 17:22:40 2024



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
