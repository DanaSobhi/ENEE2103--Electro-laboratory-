* C:\Users\CS Net Games\Desktop\4th 2ndSem\Electro lab\circuits\Prelab6N6.sch

* Schematics Version 9.1 - Web Update 1
* Sun Mar 24 18:58:40 2024



** Analysis setup **
.tran 0ns 250ms 0 10u
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Prelab6N6.net"
.INC "Prelab6N6.als"


.probe


.END
